`timescale 1ns / 1ps   // escala de tiempo [unidad de tiempo] / [precisi�n de tiempo]

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   22:17:21 09/05/2019
// Design Name:   display
// Module Name:   C:/Users/UECCI/Desktop/ejer01/display_7segx4/testbench.v
// Project Name:  display_7segx4
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: display
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module testbench;

	// Inputs
	reg [15:0] num;
	reg clk2;
	reg rst;

	// Outputs
	wire [0:6] sseg;
	wire [3:0] an;

	// Instantiate the Unit Under Test (UUT)
	display uut (  	// en este bloque llama al modulo de display y ejecuta
		.num(num), 
		.clk(clk2), 
		.sseg(sseg), 
		.an(an), 
		.rst(rst)
	);

	initial begin
		// Initialize Inputs
		clk2= 0; // apenas comienza la simulacion clk va a arrancar en cero
		rst = 1;	// apenas comienza la simulacion rst (reset) va a arrancar en uno
		#10 rst =0; //depues de un espacio de tiempo rst pasa a cero
		
		num = 16'h4321;
        

	end
      

	always #1 clk2 = ~clk2;
	
endmodule
